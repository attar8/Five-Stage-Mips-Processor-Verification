package processor_testbench_pkg;
  import uvm_pkg::*;
  
  `include "processor_sequence.sv"
  `include "processor_driver.sv"
  `include "processor_monitor.sv"
  `include "processor_scoreboard.sv"
  `include "processor_subscriber.sv"
  `include "processor_agent.sv"
  `include "processor_env.sv"
  `include "processor_test.sv"
endpackage
  
